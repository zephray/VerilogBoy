`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Wenting Zhang
// 
// Create Date:    15:28:43 02/07/2018 
// Design Name: 
// Module Name:    vga_mixer 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module vga_mixer(
    input wire clk,
    input wire rst,
    // GameBoy Image Input
    // Its clock need to be phase aligned, integer dividable by VGA clock
    // No clock domain crossing sync has been implemented here.
    input wire gb_hs,
    input wire gb_vs,
    input wire gb_pclk,
    input wire [1:0] gb_pdat,
    input wire gb_valid,
    input wire gb_en,
    // Debugger Char Input
    output wire [5:0] dbg_x,
    output wire [4:0] dbg_y,
    input wire [6:0] dbg_char,
    // VGA signal Output
    input wire pix_almost_full,
    input wire pix_next_frame,
    output wire [23:0] pix,
    output reg pix_wr,
    // Debug
    input wire hold
    );
    
    localparam GB_LIGHT = 24'h8b9a26; // Used for pixel 11
    localparam GB_MID3  = 24'h658635;
    localparam GB_MID2  = 24'h456a3e;
    localparam GB_MID1  = 24'h2d4b39;
    localparam GB_DARK  = 24'h212f25; // Used for pixel 00
    localparam GB_BACK  = 24'hbe9e16;

    //Decoded GameBoy Input colors
    wire [7:0] gb_r;
    wire [7:0] gb_g;
    wire [7:0] gb_b;
    wire [7:0] gb_grid_r;
    wire [7:0] gb_grid_g;
    wire [7:0] gb_grid_b;

    //Background colors
    wire [7:0] bg_r;
    wire [7:0] bg_g;
    wire [7:0] bg_b;

    //X,Y positions generated by the timing generator
    wire [8:0] vga_x;
    wire [8:0] vga_y;
    
    //X,Y positions of GB display
    wire [7:0] gb_x;
    wire [7:0] gb_y;

    //VGA font
    wire [6:0] font_ascii;
    wire [3:0] font_row;
    wire [2:0] font_col;
    wire font_pixel;
    
    // Font
    wire signal_in_gb_range = ((vga_y >= 16) && (vga_y < 304));
    localparam font_fg_color = 8'hFF;
    localparam font_bg_color = 8'h20;
    assign dbg_x[5:0] = vga_x[8:3];
    assign dbg_y[4:0] = vga_y[8:4];
    assign font_ascii[6:0] = dbg_char[6:0];
    assign font_row[3:0] = vga_y[3:0];
    assign font_col[2:0] = vga_x[2:0];
    wire [7:0] text_r = (font_pixel) ? (font_fg_color) : (font_bg_color);
    wire [7:0] text_g = (font_pixel) ? (font_fg_color) : (font_bg_color);
    wire [7:0] text_b = (font_pixel) ? (font_fg_color) : (font_bg_color);

    //wire is_border = (vga_x == 11'd0 || vga_x == 11'd639 || vga_y == 11'd0 || vga_y == 11'd479); 
    assign pix = (gb_en) ? ((signal_in_gb_range) ? {gb_r, gb_g, gb_b} : GB_BACK) 
            : {text_r, text_g, text_b};

    // Gameboy Input
    reg last_hold;
    
    reg [1:0] gb_buffer [0:23039];
    reg [14:0] gb_wr_addr;
    
    reg gb_vs_last;
    reg gb_hs_last;
    
    always @(posedge gb_pclk, posedge rst)
    begin
        if (rst) begin
            gb_vs_last <= 0;
            gb_hs_last <= 0;
        end
        else begin
            gb_vs_last <= gb_vs;
            gb_hs_last <= gb_hs;
        end
    end

    always @(posedge gb_pclk, posedge rst)
    begin
        if (rst) begin
            gb_wr_addr <= 0;
        end
        else begin
            if ((gb_vs_last == 1)&&(gb_vs == 0)) begin
                gb_wr_addr <= 0;
            end
            else if (gb_valid) begin
                gb_wr_addr <= gb_wr_addr + 1'b1;
                gb_buffer[gb_wr_addr] <= gb_pdat;
            end
        end
    end

    wire [14:0] gb_rd_addr = gb_y * 160 + gb_x;
    reg [1:0] gb_rd_data;
    
    always @ (posedge clk)
    begin
        gb_rd_data <= gb_buffer[gb_rd_addr];
    end
    
    assign {gb_r[7:0], gb_g[7:0], gb_b[7:0]} = 
        (gb_rd_data == 2'b11) ? (24'h212f25) : 
       ((gb_rd_data == 2'b10) ? (24'h35573e) : 
       ((gb_rd_data == 2'b01) ? (24'h597d3a) : (24'h8b9a26)));
       
    localparam X_SIZE = 320;
    localparam Y_SIZE = 320;
    
    reg [16:0] pix_counter;
    reg [8:0] x_counter;
    reg [8:0] y_counter;
    reg last_vsync;
    
    reg [7:0] red;
    reg [7:0] green;
    reg [7:0] blue;
    reg [10:0] x_raw;
    reg [9:0] x;
    
    always@(posedge clk) begin
        if (rst) begin
            pix_counter <= 0;
            pix_wr <= 1'b0;
            x_counter <= 0;
            y_counter <= 0;
        end
        else begin
            if (pix_counter < (X_SIZE * Y_SIZE)) begin
                if (pix_almost_full) begin
                    pix_wr <= 1'b0;
                end
                else begin
                    pix_counter <= pix_counter + 1;
                    if (x_counter < (X_SIZE - 1)) begin
                        x_counter <= x_counter + 1'd1;
                    end
                    else begin
                        x_counter <= 0;
                        y_counter <= y_counter + 1'd1;
                    end
                    pix_wr <= 1'b1;
                end
            end
            else begin
                pix_wr <= 1'b0;
                last_vsync <= pix_next_frame;
                if (!last_vsync && pix_next_frame) begin
                    pix_counter <= 0;
                    x_counter <= 0;
                    y_counter <= 0;
                end
            end
        end
    end
    assign vga_x = x_counter;
    assign vga_y = y_counter;
    assign gb_x = vga_x[8:1];
    assign gb_y = vga_y[8:1] - 8'd8;

    vga_font vga_font(
      .clk(clk),
      .ascii_code(font_ascii),
      .row(font_row),
      .col(font_col),
      .pixel(font_pixel)
    );    
    
endmodule
